//====================================================================
//====================== Includes ====================================
//====================================================================

//====================================================================
//============== Declaração do módulo ================================
//====================================================================

module can_crc(
	clock,
	data_in,
	enable,
	reset,
	crc
);

/** Inputs **/
input				clock;
input				data_in;
input				enable;
input				reset;

/** Outputs **/
output [14:0] crc;
reg    [14:0] crc;

/** Variáveis **/
wire          crc_next;
wire   [14:0] crc_tmp;

//====================================================================
//====================== Constantes ==================================
//====================================================================

parameter Tp = 1;

//====================================================================
//====================== Funcionamento ===============================
//====================================================================

assign crc_next = data_in ^ crc[14];
assign crc_tmp = {crc[13:0], 1'b0};

always @ (posedge clock)
begin
  if(reset)
    crc <= #Tp 15'h0;
  else if (enable)
    begin
      if (crc_next)
        crc <= #Tp crc_tmp ^ 15'h4599;
      else
        crc <= #Tp crc_tmp;
    end    
end
endmodule
