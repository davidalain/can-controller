
module bit_stuffing_framer(
	rx_bit,
	c
	tx_bit
);

input rx_bit;
output tx_bit;

wire rx_bit, tx_bit;
reg [127:0] rx_frame, [127:0] tx_frame;




endmodule
